----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    01:23:09 09/08/2022 
-- Design Name: 
-- Module Name:    Arbitro - Dataflow 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Arbitro is
	port(
		EN : in std_logic_vector(0 to 3);
		sel : out std_logic_vector(1 downto 0);
		SRC : out std_logic_vector(1 downto 0)
	);
end Arbitro;

architecture Dataflow of Arbitro is

begin
	
	sel <= "00" when EN(0) = '1' else
				"01" when EN(1) = '1' else
				"10" when EN(2) = '1' else
				"11" when EN(3) = '1';
				
	SRC <= "00" when EN(0) = '1' else
				"01" when EN(1) = '1' else
				"10" when EN(2) = '1' else
				"11" when EN(3) = '1';

end Dataflow;

